library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity TB_SecondGenerator is
end entity;

architecture behavioral of TB_SecondGenerator is

signal TB_tick_in: std_logic := '0';
signal0.