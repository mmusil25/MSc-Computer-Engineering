another_My_PLL_inst : another_My_PLL PORT MAP (
		inclk0	 => inclk0_sig,
		c0	 => c0_sig
	);
